library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fsqrttable is
  port (
    clk : in  std_logic;
    key : in  std_logic_vector(9 downto 0);
    tout : out std_logic_vector(35 downto 0) := (others => '0'));
end fsqrttable;

architecture behavioral of fsqrttable is
    type table_t is array (0 to 1023) of std_logic_vector(35 downto 0);
    constant table : table_t := (
x"6A09E969D",
x"6A6461698",
x"6ABEC1692",
x"6B190D68C",
x"6B7341687",
x"6BCD5D681",
x"6C276567C",
x"6C8155676",
x"6CDB2F671",
x"6D34F566B",
x"6D8EA1666",
x"6DE83B660",
x"6E41BD65B",
x"6E9B29655",
x"6EF481650",
x"6F4DC164A",
x"6FA6ED645",
x"700005640",
x"70590563A",
x"70B1EF635",
x"710AC5630",
x"71638562A",
x"71BC2F625",
x"7214C5620",
x"726D4561A",
x"72C5B1615",
x"731E07610",
x"73764960B",
x"73CE75605",
x"74268B600",
x"747E8D5FB",
x"74D67B5F6",
x"752E555F1",
x"7586195EB",
x"75DDC95E6",
x"7635655E1",
x"768CE95DC",
x"76E45D5D7",
x"773BBB5D2",
x"7793055CD",
x"77EA395C8",
x"7841595C3",
x"7898675BE",
x"78EF615B9",
x"7946455B4",
x"799D155AF",
x"79F3D35AA",
x"7A4A7B5A5",
x"7AA1115A0",
x"7AF79159B",
x"7B4DFF596",
x"7BA459591",
x"7BFAA158C",
x"7C50D1587",
x"7CA6F1582",
x"7CFCFD57E",
x"7D52F5579",
x"7DA8DB574",
x"7DFEAD56F",
x"7E546B56A",
x"7EAA15566",
x"7EFFAD561",
x"7F553355C",
x"7FAAA5557",
x"800003552",
x"80554F54E",
x"80AA89549",
x"80FFAD544",
x"8154C1540",
x"81A9C153B",
x"81FEB1536",
x"82538B532",
x"82A85352D",
x"82FD09528",
x"8351AD524",
x"83A63D51F",
x"83FABD51B",
x"844F29516",
x"84A381511",
x"84F7C950D",
x"854BFD508",
x"85A021504",
x"85F4314FF",
x"8648314FB",
x"869C1D4F6",
x"86EFF94F2",
x"8743C14ED",
x"8797794E9",
x"87EB1D4E4",
x"883EB14E0",
x"8892314DB",
x"88E5A14D7",
x"8938FD4D3",
x"898C4B4CE",
x"89DF854CA",
x"8A32AD4C5",
x"8A85C54C1",
x"8AD8CB4BD",
x"8B2BC14B8",
x"8B7EA34B4",
x"8BD1754B0",
x"8C24354AB",
x"8C76E54A7",
x"8CC9814A3",
x"8D1C0F49E",
x"8D6E8B49A",
x"8DC0F5496",
x"8E134F492",
x"8E659748D",
x"8EB7CD489",
x"8F09F5485",
x"8F5C09481",
x"8FAE0F47C",
x"900003478",
x"9051E5474",
x"90A3B9470",
x"90F57946C",
x"91472B468",
x"9198CD463",
x"91EA5D45F",
x"923BDB45B",
x"928D49457",
x"92DEA9453",
x"932FF544F",
x"93813544B",
x"93D261447",
x"94237D443",
x"94748943F",
x"94C58743B",
x"951673437",
x"95674F432",
x"95B81B42E",
x"9608D742A",
x"965983426",
x"96AA1D422",
x"96FAA941E",
x"974B2541B",
x"979B91417",
x"97EBED413",
x"983C3B40F",
x"988C7740B",
x"98DCA5407",
x"992CC1403",
x"997CCF3FF",
x"99CCCD3FB",
x"9A1CBB3F7",
x"9A6C993F3",
x"9ABC693EF",
x"9B0C293EC",
x"9B5BD93E8",
x"9BAB793E4",
x"9BFB093E0",
x"9C4A8D3DC",
x"9C99FF3D8",
x"9CE9613D5",
x"9D38B53D1",
x"9D87FB3CD",
x"9DD7313C9",
x"9E26593C5",
x"9E756F3C2",
x"9EC4793BE",
x"9F13713BA",
x"9F625B3B6",
x"9FB1353B3",
x"A000033AF",
x"A04EC13AB",
x"A09D6F3A7",
x"A0EC0F3A4",
x"A13AA13A0",
x"A1892139C",
x"A1D795399",
x"A225F9395",
x"A27451391",
x"A2C29738E",
x"A310D138A",
x"A35EF9386",
x"A3AD15383",
x"A3FB2137F",
x"A4492137C",
x"A49711378",
x"A4E4F3374",
x"A532C5371",
x"A5808B36D",
x"A5CE4136A",
x"A61BE9366",
x"A66985362",
x"A6B70F35F",
x"A7048D35B",
x"A751FD358",
x"A79F5D354",
x"A7ECB1351",
x"A839F534D",
x"A8872D34A",
x"A8D455346",
x"A92171343",
x"A96E7D33F",
x"A9BB7B33C",
x"AA086D338",
x"AA5551335",
x"AAA225331",
x"AAEEED32E",
x"AB3BA532A",
x"AB8851327",
x"ABD4F1324",
x"AC2181320",
x"AC6E0331D",
x"ACBA79319",
x"AD06DF316",
x"AD5339313",
x"AD9F8530F",
x"ADEBC530C",
x"AE37F5308",
x"AE8419305",
x"AED031302",
x"AF1C392FE",
x"AF68352FB",
x"AFB4212F8",
x"B000032F4",
x"B04BD52F1",
x"B0979D2EE",
x"B0E3552EA",
x"B12F012E7",
x"B17A9F2E4",
x"B1C6312E1",
x"B211B52DD",
x"B25D2B2DA",
x"B2A8952D7",
x"B2F3F12D3",
x"B33F412D0",
x"B38A852CD",
x"B3D5B92CA",
x"B420E32C6",
x"B46BFF2C3",
x"B4B70D2C0",
x"B5020F2BD",
x"B54D052BA",
x"B597ED2B6",
x"B5E2C92B3",
x"B62D972B0",
x"B678592AD",
x"B6C30D2AA",
x"B70DB72A6",
x"B758512A3",
x"B7A2E12A0",
x"B7ED6529D",
x"B837D929A",
x"B88243297",
x"B8CCA1294",
x"B916F1290",
x"B9613528D",
x"B9AB6B28A",
x"B9F595287",
x"BA3FB5284",
x"BA89C5281",
x"BAD3CB27E",
x"BB1DC527B",
x"BB67B1278",
x"BBB191275",
x"BBFB65271",
x"BC452D26E",
x"BC8EE926B",
x"BCD899268",
x"BD223D265",
x"BD6BD3262",
x"BDB55D25F",
x"BDFEDD25C",
x"BE484F259",
x"BE91B5256",
x"BEDB11253",
x"BF245F250",
x"BF6DA124D",
x"BFB6D924A",
x"C00001247",
x"C04921244",
x"C09235241",
x"C0DB3B23E",
x"C1243523B",
x"C16D25238",
x"C1B609235",
x"C1FEDF232",
x"C247AB22F",
x"C2906B22D",
x"C2D91F22A",
x"C321C7227",
x"C36A65224",
x"C3B2F5221",
x"C3FB7B21E",
x"C443F521B",
x"C48C61218",
x"C4D4C5215",
x"C51D1D212",
x"C5656920F",
x"C5ADA920D",
x"C5F5DD20A",
x"C63E05207",
x"C68621204",
x"C6CE35201",
x"C7163B1FE",
x"C75E371FB",
x"C7A6251F9",
x"C7EE0B1F6",
x"C835E51F3",
x"C87DB11F0",
x"C8C5751ED",
x"C90D2D1EB",
x"C954D91E8",
x"C99C791E5",
x"C9E40F1E2",
x"CA2B991DF",
x"CA73191DD",
x"CABA8D1DA",
x"CB01F51D7",
x"CB49551D4",
x"CB90A71D1",
x"CBD7EF1CF",
x"CC1F2D1CC",
x"CC665D1C9",
x"CCAD851C6",
x"CCF4A11C4",
x"CD3BB11C1",
x"CD82B71BE",
x"CDC9B11BC",
x"CE10A11B9",
x"CE57871B6",
x"CE9E611B3",
x"CEE5311B1",
x"CF2BF51AE",
x"CF72AF1AB",
x"CFB95D1A9",
x"D000011A6",
x"D0469D1A3",
x"D08D2B1A1",
x"D0D3AF19E",
x"D11A2919B",
x"D16097199",
x"D1A6FB196",
x"D1ED55193",
x"D233A3191",
x"D279E718E",
x"D2C02118B",
x"D30651189",
x"D34C75186",
x"D3928F183",
x"D3D89D181",
x"D41EA317E",
x"D4649D17C",
x"D4AA8D179",
x"D4F075176",
x"D5364F174",
x"D57C21171",
x"D5C1E516F",
x"D607A116C",
x"D64D55169",
x"D692FD167",
x"D6D899164",
x"D71E2D162",
x"D763B515F",
x"D7A93315D",
x"D7EEA715A",
x"D83411157",
x"D87971155",
x"D8BEC5152",
x"D90411150",
x"D9495314D",
x"D98E8914B",
x"D9D3B7148",
x"DA18D9146",
x"DA5DF1143",
x"DAA301141",
x"DAE80513E",
x"DB2D0113C",
x"DB71F1139",
x"DBB6D9137",
x"DBFBB5134",
x"DC4089132",
x"DC855112F",
x"DCCA0F12D",
x"DD0EC512A",
x"DD536F128",
x"DD9811125",
x"DDDCA9123",
x"DE2135120",
x"DE65B911E",
x"DEAA3311C",
x"DEEEA3119",
x"DF3309117",
x"DF7765114",
x"DFBBB9112",
x"E0000110F",
x"E0444110D",
x"E0887710B",
x"E0CCA3108",
x"E110C5106",
x"E154DF103",
x"E198ED101",
x"E1DCF30FE",
x"E220EF0FC",
x"E264E10FA",
x"E2A8C90F7",
x"E2ECA90F5",
x"E3307F0F3",
x"E3744B0F0",
x"E3B80D0EE",
x"E3FBC70EB",
x"E43F770E9",
x"E4831D0E7",
x"E4C6B90E4",
x"E50A4D0E2",
x"E54DD70E0",
x"E591590DD",
x"E5D4CF0DB",
x"E6183D0D9",
x"E65BA10D6",
x"E69EFD0D4",
x"E6E24D0D2",
x"E725970CF",
x"E768D50CD",
x"E7AC0D0CB",
x"E7EF390C8",
x"E8325D0C6",
x"E875750C4",
x"E8B8870C1",
x"E8FB8F0BF",
x"E93E8D0BD",
x"E981830BB",
x"E9C46F0B8",
x"EA07530B6",
x"EA4A2D0B4",
x"EA8CFD0B1",
x"EACFC50AF",
x"EB12850AD",
x"EB55390AB",
x"EB97E50A8",
x"EBDA890A6",
x"EC1D250A4",
x"EC5FB50A2",
x"ECA23F09F",
x"ECE4BD09D",
x"ED273509B",
x"ED69A3099",
x"EDAC07096",
x"EDEE63094",
x"EE30B5092",
x"EE7301090",
x"EEB54108E",
x"EEF77908B",
x"EF39A9089",
x"EF7BCF087",
x"EFBDED085",
x"F00001083",
x"F0420D080",
x"F0841107E",
x"F0C60D07C",
x"F107FD07A",
x"F149E7078",
x"F18BC7075",
x"F1CD9F073",
x"F20F6D071",
x"F2513506F",
x"F292F106D",
x"F2D4A506B",
x"F31653068",
x"F357F5066",
x"F39991064",
x"F3DB25062",
x"F41CAD060",
x"F45E2D05E",
x"F49FA705C",
x"F4E117059",
x"F5227F057",
x"F563DD055",
x"F5A535053",
x"F5E681051",
x"F627C704F",
x"F6690504D",
x"F6AA3904B",
x"F6EB65048",
x"F72C89046",
x"F76DA5044",
x"F7AEB5042",
x"F7EFC1040",
x"F830C303E",
x"F871BD03C",
x"F8B2AD03A",
x"F8F395038",
x"F93477036",
x"F9754F033",
x"F9B61F031",
x"F9F6E702F",
x"FA37A502D",
x"FA785D02B",
x"FAB90D029",
x"FAF9B1027",
x"FB3A51025",
x"FB7AE7023",
x"FBBB75021",
x"FBFBF901F",
x"FC3C7701D",
x"FC7CED01B",
x"FCBD59019",
x"FCFDBF017",
x"FD3E1B015",
x"FD7E71013",
x"FDBEBD011",
x"FDFF0100F",
x"FE3F3D00D",
x"FE7F7100B",
x"FEBF9D009",
x"FEFFC1007",
x"FF3FDD005",
x"FF7FF1003",
x"FFBFFD001",
x"000002FFE",
x"003FFAFFA",
x"007FE2FF6",
x"00BFBAFF2",
x"00FF82FEE",
x"013F3CFEA",
x"017EE4FE6",
x"01BE7CFE2",
x"01FE06FDE",
x"023D80FDA",
x"027CEAFD6",
x"02BC44FD2",
x"02FB90FCE",
x"033ACCFCB",
x"0379F8FC7",
x"03B914FC3",
x"03F820FBF",
x"043720FBB",
x"04760EFB7",
x"04B4EEFB4",
x"04F3C0FB0",
x"053280FAC",
x"057134FA8",
x"05AFD6FA5",
x"05EE6CFA1",
x"062CF0F9D",
x"066B68F99",
x"06A9D0F96",
x"06E828F92",
x"072672F8E",
x"0764ACF8B",
x"07A2DAF87",
x"07E0F8F83",
x"081F08F80",
x"085D08F7C",
x"089AFCF78",
x"08D8E0F75",
x"0916B4F71",
x"09547CF6E",
x"099234F6A",
x"09CFE0F67",
x"0A0D7CF63",
x"0A4B08F5F",
x"0A8888F5C",
x"0AC5FAF58",
x"0B035CF55",
x"0B40B2F51",
x"0B7DF8F4E",
x"0BBB32F4A",
x"0BF85CF47",
x"0C357AF43",
x"0C728AF40",
x"0CAF8CF3C",
x"0CEC80F39",
x"0D2964F35",
x"0D663CF32",
x"0DA308F2F",
x"0DDFC4F2B",
x"0E1C72F28",
x"0E5914F24",
x"0E95A8F21",
x"0ED22CF1E",
x"0F0EA6F1A",
x"0F4B10F17",
x"0F876EF14",
x"0FC3C0F10",
x"100002F0D",
x"103C38F0A",
x"107860F06",
x"10B47AF03",
x"10F088F00",
x"112C88EFC",
x"11687CEF9",
x"11A462EF6",
x"11E03CEF3",
x"121C08EEF",
x"1257C8EEC",
x"129378EE9",
x"12CF1EEE6",
x"130AB6EE2",
x"134640EDF",
x"1381C0EDC",
x"13BD30ED9",
x"13F896ED5",
x"1433EEED2",
x"146F38ECF",
x"14AA78ECC",
x"14E5A8EC9",
x"1520D0EC6",
x"155BE8EC3",
x"1596F4EBF",
x"15D1F4EBC",
x"160CE6EB9",
x"1647CCEB6",
x"1682A6EB3",
x"16BD74EB0",
x"16F834EAD",
x"1732EAEAA",
x"176D92EA7",
x"17A82EEA3",
x"17E2BEEA0",
x"181D42E9D",
x"1857B8E9A",
x"189224E97",
x"18CC84E94",
x"1906D8E91",
x"19411CE8E",
x"197B58E8B",
x"19B588E88",
x"19EFAAE85",
x"1A29C0E82",
x"1A63CCE7F",
x"1A9DCAE7C",
x"1AD7BCE79",
x"1B11A4E76",
x"1B4B80E73",
x"1B8550E70",
x"1BBF14E6E",
x"1BF8CCE6B",
x"1C3278E68",
x"1C6C18E65",
x"1CA5ACE62",
x"1CDF36E5F",
x"1D18B4E5C",
x"1D5226E59",
x"1D8B8CE56",
x"1DC4E8E53",
x"1DFE38E51",
x"1E377CE4E",
x"1E70B4E4B",
x"1EA9E0E48",
x"1EE304E45",
x"1F1C18E42",
x"1F5524E3F",
x"1F8E24E3D",
x"1FC718E3A",
x"200000E37",
x"2038E0E34",
x"2071B2E31",
x"20AA7AE2F",
x"20E336E2C",
x"211BE8E29",
x"21548CE26",
x"218D28E24",
x"21C5B8E21",
x"21FE3CE1E",
x"2236B8E1B",
x"226F26E19",
x"22A78AE16",
x"22DFE4E13",
x"231832E10",
x"235074E0E",
x"2388ACE0B",
x"23C0DCE08",
x"23F8FEE06",
x"243116E03",
x"246924E00",
x"24A126DFD",
x"24D91CDFB",
x"25110ADF8",
x"2548ECDF5",
x"2580C4DF3",
x"25B892DF0",
x"25F054DEE",
x"26280CDEB",
x"265FBADE8",
x"26975CDE6",
x"26CEF4DE3",
x"270684DE0",
x"273E08DDE",
x"277580DDB",
x"27ACF0DD9",
x"27E454DD6",
x"281BACDD3",
x"2852FCDD1",
x"288A42DCE",
x"28C17CDCC",
x"28F8AEDC9",
x"292FD4DC7",
x"2966F0DC4",
x"299E02DC1",
x"29D50ADBF",
x"2A0C08DBC",
x"2A42FCDBA",
x"2A79E4DB7",
x"2AB0C4DB5",
x"2AE79ADB2",
x"2B1E64DB0",
x"2B5526DAD",
x"2B8BDCDAB",
x"2BC28ADA8",
x"2BF92EDA6",
x"2C2FC8DA3",
x"2C6656DA1",
x"2C9CDCD9E",
x"2CD358D9C",
x"2D09C8D99",
x"2D4030D97",
x"2D7690D95",
x"2DACE4D92",
x"2DE32ED90",
x"2E196ED8D",
x"2E4FA4D8B",
x"2E85D4D88",
x"2EBBF6D86",
x"2EF210D84",
x"2F2820D81",
x"2F5E28D7F",
x"2F9424D7C",
x"2FCA18D7A",
x"300000D78",
x"3035E0D75",
x"306BB8D73",
x"30A184D70",
x"30D748D6E",
x"310D04D6C",
x"3142B4D69",
x"31785CD67",
x"31ADFAD65",
x"31E38ED62",
x"321918D60",
x"324E9CD5E",
x"328414D5B",
x"32B984D59",
x"32EEE8D57",
x"332444D54",
x"335998D52",
x"338EE2D50",
x"33C424D4D",
x"33F95CD4B",
x"342E88D49",
x"3463B0D47",
x"3498CCD44",
x"34CDDED42",
x"3502E8D40",
x"3537E8D3D",
x"356CE0D3B",
x"35A1CED39",
x"35D6B4D37",
x"360B90D34",
x"364064D32",
x"367530D30",
x"36A9F0D2E",
x"36DEA8D2B",
x"371358D29",
x"374800D27",
x"377C9CD25",
x"37B132D23",
x"37E5BED20",
x"381A42D1E",
x"384EBCD1C",
x"38832ED1A",
x"38B798D18",
x"38EBF8D15",
x"39204ED13",
x"39549CD11",
x"3988E2D0F",
x"39BD20D0D",
x"39F154D0A",
x"3A2580D08",
x"3A59A4D06",
x"3A8DBCD04",
x"3AC1D0D02",
x"3AF5D8D00",
x"3B29D8CFE",
x"3B5DD0CFB",
x"3B91C0CF9",
x"3BC5A8CF7",
x"3BF986CF5",
x"3C2D5CCF3",
x"3C6128CF1",
x"3C94EECEF",
x"3CC8ACCED",
x"3CFC60CEA",
x"3D300ACE8",
x"3D63AECE6",
x"3D9748CE4",
x"3DCADCCE2",
x"3DFE64CE0",
x"3E31E8CDE",
x"3E6560CDC",
x"3E98D0CDA",
x"3ECC3ACD8",
x"3EFF9ACD6",
x"3F32F4CD3",
x"3F6642CD1",
x"3F998ACCF",
x"3FCCCACCD",
x"400000CCB",
x"403330CC9",
x"406658CC7",
x"409976CC5",
x"40CC8CCC3",
x"40FF9CCC1",
x"4132A0CBF",
x"4165A0CBD",
x"419896CBB",
x"41CB84CB9",
x"41FE6ACB7",
x"423148CB5",
x"42641ECB3",
x"4296ECCB1",
x"42C9B2CAF",
x"42FC70CAD",
x"432F26CAB",
x"4361D4CA9",
x"43947ACA7",
x"43C718CA5",
x"43F9B0CA3",
x"442C3CCA1",
x"445EC4C9F",
x"449142C9D",
x"44C3B8C9B",
x"44F628C99",
x"452890C97",
x"455AF0C95",
x"458D46C93",
x"45BF96C92",
x"45F1DEC90",
x"46241EC8E",
x"465658C8C",
x"468888C8A",
x"46BAB0C88",
x"46ECD2C86",
x"471EECC84",
x"4750FEC82",
x"478308C80",
x"47B50CC7E",
x"47E706C7C",
x"4818FAC7A",
x"484AE6C79",
x"487CCAC77",
x"48AEA8C75",
x"48E07CC73",
x"49124AC71",
x"494410C6F",
x"4975CEC6D",
x"49A784C6B",
x"49D934C6A",
x"4A0ADCC68",
x"4A3C7EC66",
x"4A6E18C64",
x"4A9FA8C62",
x"4AD134C60",
x"4B02B6C5E",
x"4B3430C5D",
x"4B65A6C5B",
x"4B9712C59",
x"4BC878C57",
x"4BF9D6C55",
x"4C2B2CC53",
x"4C5C7CC52",
x"4C8DC4C50",
x"4CBF04C4E",
x"4CF03EC4C",
x"4D2170C4A",
x"4D529CC48",
x"4D83C0C47",
x"4DB4DCC45",
x"4DE5F0C43",
x"4E1700C41",
x"4E4804C3F",
x"4E7904C3E",
x"4EA9FCC3C",
x"4EDAF0C3A",
x"4F0BD8C38",
x"4F3CBCC36",
x"4F6D98C35",
x"4F9E6CC33",
x"4FCF3AC31",
x"500000C2F",
x"5030C0C2E",
x"506178C2C",
x"50922AC2A",
x"50C2D4C28",
x"50F378C27",
x"512414C25",
x"5154AAC23",
x"518538C21",
x"51B5C0C20",
x"51E640C1E",
x"5216B8C1C",
x"52472CC1A",
x"527798C19",
x"52A7FCC17",
x"52D858C15",
x"5308B0C13",
x"533900C12",
x"536948C10",
x"53998CC0E",
x"53C9C6C0D",
x"53F9FCC0B",
x"542A28C09",
x"545A50C08",
x"548A70C06",
x"54BA88C04",
x"54EA9CC02",
x"551AA6C01",
x"554AACBFF",
x"557AA8BFD",
x"55AAA0BFC",
x"55DA92BFA",
x"560A7CBF8",
x"563A60BF7",
x"566A3CBF5",
x"569A10BF3",
x"56C9E0BF2",
x"56F9A8BF0",
x"57296CBEE",
x"575926BED",
x"5788DABEB",
x"57B888BE9",
x"57E830BE8",
x"5817D0BE6",
x"58476CBE4",
x"5876FEBE3",
x"58A68CBE1",
x"58D612BDF",
x"590590BDE",
x"59350CBDC",
x"59647EBDB",
x"5993EABD9",
x"59C350BD7",
x"59F2B0BD6",
x"5A2208BD4",
x"5A515ABD2",
x"5A80A6BD1",
x"5AAFECBCF",
x"5ADF2CBCE",
x"5B0E64BCC",
x"5B3D96BCA",
x"5B6CC0BC9",
x"5B9BE8BC7",
x"5BCB06BC6",
x"5BFA1EBC4",
x"5C2930BC2",
x"5C583CBC1",
x"5C8742BBF",
x"5CB640BBE",
x"5CE53ABBC",
x"5D142CBBB",
x"5D4318BB9",
x"5D71FEBB7",
x"5DA0DEBB6",
x"5DCFB8BB4",
x"5DFE8ABB3",
x"5E2D58BB1",
x"5E5C1EBB0",
x"5E8ADEBAE",
x"5EB998BAC",
x"5EE84CBAB",
x"5F16F8BA9",
x"5F45A0BA8",
x"5F7442BA6",
x"5FA2DCBA5",
x"5FD172BA3",
x"600000BA2",
x"602E88BA0",
x"605D0CB9F",
x"608B88B9D",
x"60B9FEB9C",
x"60E86EB9A",
x"6116D8B98",
x"61453CB97",
x"61739AB95",
x"61A1F0B94",
x"61D044B92",
x"61FE8EB91",
x"622CD4B8F",
x"625B14B8E",
x"62894CB8C",
x"62B780B8B",
x"62E5AEB89",
x"6313D4B88",
x"6341F6B86",
x"637012B85",
x"639E28B83",
x"63CC38B82",
x"63FA40B80",
x"642844B7F",
x"645640B7D",
x"648438B7C",
x"64B22AB7A",
x"64E016B79",
x"650DFCB78",
x"653BDCB76",
x"6569B6B75",
x"65978CB73",
x"65C558B72",
x"65F320B70",
x"6620E4B6F",
x"664EA0B6D",
x"667C58B6C",
x"66AA08B6A",
x"66D7B4B69",
x"67055AB67",
x"6732FAB66",
x"676094B65",
x"678E28B63",
x"67BBB6B62",
x"67E940B60",
x"6816C0B5F",
x"684440B5D",
x"6871B6B5C",
x"689F28B5A",
x"68CC94B59",
x"68F9FAB58",
x"69275AB56",
x"6954B4B55",
x"69820AB53",
x"69AF58B52",
x"69DCA4B51");

begin
    process(key)
    begin
       -- if rising_edge(clk) then
            tout <= table(to_integer(unsigned(key)));
       -- end if;
    end process;
end behavioral;
